package Cafe;

// The only argument to the cafe function is the size of t.
import "BDPI" cafe = function ActionValue#(t) cafe_c (Bit#(32) sz)
  provisos (Bits#(t, sz));

endpackage