package Beef;

// The only argument to the beef function is the size of t.
import "BDPI" beef = function ActionValue#(t) beef_c (Bit#(32) sz)
  provisos (Bits#(t, sz));

endpackage