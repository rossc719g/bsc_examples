package Raw where

data Raw t = Raw (Bit (SizeOf t))

instance (Bits t sz) => Bits (Raw t) sz where
  pack   (Raw x) = x
  unpack x       = Raw x

instance (Bits t tsz) => DefaultValue (Raw t) where
  defaultValue = Raw defaultValue

cook :: (Bits t tsz) => Raw t -> t
cook (Raw x) = unpack x

uncook :: (Bits t tsz) => t -> Raw t
uncook x = Raw (pack x)
